
# run -all
# time=0| tx_start=0 | tx_data=0| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=idle 
# time=104170| tx_start=1 | tx_data=36| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=idle 
# time=104190| tx_start=0 | tx_data=36| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=start 
# time=208350| tx_start=0 | tx_data=36| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=data 
# time=416670| tx_start=0 | tx_data=36| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=data 
# time=520830| tx_start=0 | tx_data=36| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=data 
# time=729150| tx_start=0 | tx_data=36| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=data 
# time=833310| tx_start=0 | tx_data=36| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=data 
# time=1041630| tx_start=0 | tx_data=36| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=parity 
# time=1145790| tx_start=0 | tx_data=36| tx_out=1| tx_done=1| rx_done=0| rx_data_out=(  x)xxxxxxxx |tx_state=stop 
# time=1196030| tx_start=0 | tx_data=36| tx_out=1| tx_done=1| rx_done=1| rx_data_out=(  x)xxxxxxxx |tx_state=stop 
# time=1196050| tx_start=0 | tx_data=36| tx_out=1| tx_done=1| rx_done=1| rx_data_out=( 36)00100100 |tx_state=stop 
# time=1202530| tx_start=0 | tx_data=36| tx_out=1| tx_done=1| rx_done=0| rx_data_out=( 36)00100100 |tx_state=stop 
# time=1249930| tx_start=1 | tx_data=1| tx_out=1| tx_done=1| rx_done=0| rx_data_out=( 36)00100100 |tx_state=stop 

# time=1249950| tx_start=0 | tx_data=1| tx_out=0| tx_done=0| rx_done=0| rx_data_out=( 36)00100100 |tx_state=start 
# time=1354110| tx_start=0 | tx_data=1| tx_out=1| tx_done=0| rx_done=0| rx_data_out=( 36)00100100 |tx_state=data 
# time=1458270| tx_start=0 | tx_data=1| tx_out=0| tx_done=0| rx_done=0| rx_data_out=( 36)00100100 |tx_state=data 
# time=2187390| tx_start=0 | tx_data=1| tx_out=1| tx_done=0| rx_done=0| rx_data_out=( 36)00100100 |tx_state=parity 
# time=2291550| tx_start=0 | tx_data=1| tx_out=1| tx_done=1| rx_done=0| rx_data_out=( 36)00100100 |tx_state=stop 
# time=2340030| tx_start=0 | tx_data=1| tx_out=1| tx_done=1| rx_done=1| rx_data_out=( 36)00100100 |tx_state=stop 
# time=2340050| tx_start=0 | tx_data=1| tx_out=1| tx_done=1| rx_done=1| rx_data_out=(  1)00000001 |tx_state=stop 
# time=2346530| tx_start=0 | tx_data=1| tx_out=1| tx_done=1| rx_done=0| rx_data_out=(  1)00000001 |tx_state=stop 
# time=2395690| tx_start=1 | tx_data=9| tx_out=1| tx_done=1| rx_done=0| rx_data_out=(  1)00000001 |tx_state=stop 

# time=2395710| tx_start=0 | tx_data=9| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=start 
# time=2499870| tx_start=0 | tx_data=9| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=data 
# time=2604030| tx_start=0 | tx_data=9| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=data 
# time=2812350| tx_start=0 | tx_data=9| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=data 
# time=2916510| tx_start=0 | tx_data=9| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=data 
# time=3333150| tx_start=0 | tx_data=9| tx_out=0| tx_done=0| rx_done=0| rx_data_out=(  1)00000001 |tx_state=parity 
# time=3437310| tx_start=0 | tx_data=9| tx_out=1| tx_done=1| rx_done=0| rx_data_out=(  1)00000001 |tx_state=stop 
# time=3484030| tx_start=0 | tx_data=9| tx_out=1| tx_done=1| rx_done=1| rx_data_out=(  1)00000001 |tx_state=stop 
# time=3484050| tx_start=0 | tx_data=9| tx_out=1| tx_done=1| rx_done=1| rx_data_out=(  9)00001001 |tx_state=stop 
# time=3490530| tx_start=0 | tx_data=9| tx_out=1| tx_done=1| rx_done=0| rx_data_out=(  9)00001001 |tx_state=stop 
# time=3541470| tx_start=0 | tx_data=9| tx_out=1| tx_done=0| rx_done=0| rx_data_out=(  9)00001001 |tx_state=idle 
# ** Note: $finish    : testbench.sv(53)
#    Time: 5437310 ns  Iteration: 0  Instance: /uart_tb
